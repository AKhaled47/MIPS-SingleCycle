module instruction_mem(
    input [31:0] Address,
    output [31:0] RD
);

wire [5:0] shifted_address;
assign shifted_address = Address [7:2];
wire [31:0] INS_MEM [0:44];




assign INS_MEM[0] = 32'b00100000000010000000000000010000; //Begin:  addi t0 zero 0x10    16
assign INS_MEM[1] = 32'b00100000000010010000000000001010; //        addi t1 zero 0x0a    10
assign INS_MEM[2] = 32'b00000001000010011000000000100100; //        and $s0, $t0, $t1    0
assign INS_MEM[3] = 32'b00000001000010011000000000100101; //        or $s0, $t0, $t1    26
assign INS_MEM[4] = 32'b10101100000100000000000000000100; //        sw $s0, 4($zero)  4  
assign INS_MEM[5] = 32'b10101100000010000000000000001000; //        sw $t0, 8($zero)    8
assign INS_MEM[6] = 32'b00000001000010011000100000100000; //        add $s1, $t0, $t1    26 
assign INS_MEM[7] = 32'b00000001000010011001000000100010; //        sub $s2, $t0, $t1    6
assign INS_MEM[8] = 32'b10001100000100010000000000000100; //        lw $s1, 4($zero)    26
assign INS_MEM[9] = 32'b00100010001100100000000001001000; //        addi $s2, $s1, 0x48   98  
assign INS_MEM[10] = 32'b10001100000100110000000000001000; //       lw $s3, 8($zero)    16
assign INS_MEM[11] = 32'b00000010001100111001000000100000; //       add s2 s1 s3     42
assign INS_MEM[12] = 32'b00000000000000001000100000100000 ;//       add $s1 $0 $0    0
assign INS_MEM[13] = 32'b00000000000000001000000000100000 ;//       add $s0 $0 $0     0
assign INS_MEM[14] = 32'b00100000000010000000000000001010; //       add $t0 $0 $10     0
assign INS_MEM[15] = 32'b00010001000100000000000000000011; //for:   beq $s0, $t0, done                         
assign INS_MEM[16] = 32'b00000010001100001000100000100000 ;//       add $s1 $s1 $s0          
assign INS_MEM[17] = 32'b00100010000100000000000000000001 ;//       ADDI $s0 $s0 0x1                                            
assign INS_MEM[18] = 32'b00001000000000000000000000001111 ; //      j for  
assign INS_MEM[19] = 32'b00001000000000000000000000000000; //done : j Begin              



//********************************************************************************************************************************

/*


assign INS_MEM[0] = 32'b00100000000010010000000000001111; //addi t1 zero 0x0f    15
assign INS_MEM[1] = 32'b00000000000000001000100000100000 ;//add $s1 $0 $0    0
assign INS_MEM[2] = 32'b00000000000000001000000000100000 ;//add $s0 $0 $0     0
assign INS_MEM[3] = 32'b00100000000010000000000000001010; //add $t0 $0 $10     0
assign INS_MEM[4] = 32'b00010001000100000000000000000011;    //for:     beq $s0, $t0, done                         
assign INS_MEM[5] = 32'b00000010001100001000100000100000 ;//add $s1 $s1 $s0          
assign INS_MEM[6] = 32'b00100010000100000000000000000001 ;//ADDI $s0 $s0 0x1                                            
assign INS_MEM[7] = 32'b00001000000000000000000000000100; //j for  
assign INS_MEM[8] = 32'b00001000000000000000000000000000; //j Begin                      
*/





//******************************************************************************************



assign RD = INS_MEM [shifted_address];

endmodule